module node_op(
  input logic  clk,
  input logic  rst,
  input logic valid_in,

  input logic prev_outputs,
  input logic weigths,
  input logic biases,
  
  output logic valid_out,
  output logic x,
);


  // load all (3?) arrays
  //do first calculation and load
  //dp second calculation and load

  
